library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package util_package is    
    function sbox (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function T (j:integer;x:std_logic_vector(31 downto 0)) return std_logic_vector;
end util_package;

package body util_package is
-------------transform function for key expansion---------
function T (j:integer;x:std_logic_vector(31 downto 0)) return std_logic_vector is
    variable a:std_logic_vector(31 downto 0);
    variable b:std_logic_vector(31 downto 0);
    variable c:std_logic_vector(31 downto 0);
begin
    a:=x(23 downto 0)&x(31 downto 24);
    b:=sbox(a(31 downto 24)) & sbox(a(23 downto 16)) & sbox(a(15 downto 8)) & sbox(a(7 downto 0));
    case j is
        when 1 => c:= "00000001000000000000000000000000" xor b;
        when 2 => c:= "00000010000000000000000000000000" xor b;
        when 3 => c:= "00000100000000000000000000000000" xor b;
        when 4 => c:= "00001000000000000000000000000000" xor b;
        when 5 => c:= "00010000000000000000000000000000" xor b;
        when 6 => c:= "00100000000000000000000000000000" xor b;
        when 7 => c:= "01000000000000000000000000000000" xor b;
        when 8 => c:= "10000000000000000000000000000000" xor b;
        when 9 => c:= "00011011000000000000000000000000" xor b;
        when 10=> c:= "00110110000000000000000000000000" xor b;
        when others => c:="00000000000000000000000000000000";
    end case;
    return c;
end function;

-----------sbox function (created for functions above)------
function sbox (x: std_logic_vector(7 downto 0)) return std_logic_vector is 
    variable i:std_logic_vector(7 downto 0);
begin
    case x is
        when x"00" =>i:=x"63";
		when x"01" =>i:=x"7c";
		when x"02" =>i:=x"77";
		when x"03" =>i:=x"7b";
		when x"04" =>i:=x"f2";
		when x"05" =>i:=x"6b";
		when x"06" =>i:=x"6f";
		when x"07" =>i:=x"c5";
		when x"08" =>i:=x"30";
		when x"09" =>i:=x"01";
		when x"0a" =>i:=x"67";
		when x"0b" =>i:=x"2b";
		when x"0c" =>i:=x"fe";
		when x"0d" =>i:=x"d7";
		when x"0e" =>i:=x"ab";
		when x"0f" =>i:=x"76";
		when x"10" =>i:=x"ca";
		when x"11" =>i:=x"82";
		when x"12" =>i:=x"c9";
		when x"13" =>i:=x"7d";
		when x"14" =>i:=x"fa";
		when x"15" =>i:=x"59";
		when x"16" =>i:=x"47";
		when x"17" =>i:=x"f0";
		when x"18" =>i:=x"ad";
		when x"19" =>i:=x"d4";
		when x"1a" =>i:=x"a2";
		when x"1b" =>i:=x"af";
		when x"1c" =>i:=x"9c";
		when x"1d" =>i:=x"a4";
		when x"1e" =>i:=x"72";
		when x"1f" =>i:=x"c0";
		when x"20" =>i:=x"b7";
		when x"21" =>i:=x"fd";
		when x"22" =>i:=x"93";
		when x"23" =>i:=x"26";
		when x"24" =>i:=x"36";
		when x"25" =>i:=x"3f";
		when x"26" =>i:=x"f7";
		when x"27" =>i:=x"cc";
		when x"28" =>i:=x"34";
		when x"29" =>i:=x"a5";
		when x"2a" =>i:=x"e5";
		when x"2b" =>i:=x"f1";
		when x"2c" =>i:=x"71";
		when x"2d" =>i:=x"d8";
		when x"2e" =>i:=x"31";
		when x"2f" =>i:=x"15";
		when x"30" =>i:=x"04";
		when x"31" =>i:=x"c7";
		when x"32" =>i:=x"23";
		when x"33" =>i:=x"c3";
		when x"34" =>i:=x"18";
		when x"35" =>i:=x"96";
		when x"36" =>i:=x"05";
		when x"37" =>i:=x"9a";
		when x"38" =>i:=x"07";
		when x"39" =>i:=x"12";
		when x"3a" =>i:=x"80";
		when x"3b" =>i:=x"e2";
		when x"3c" =>i:=x"eb";
		when x"3d" =>i:=x"27";
		when x"3e" =>i:=x"b2";
		when x"3f" =>i:=x"75";
		when x"40" =>i:=x"09";
		when x"41" =>i:=x"83";
		when x"42" =>i:=x"2c";
		when x"43" =>i:=x"1a";
		when x"44" =>i:=x"1b";
		when x"45" =>i:=x"6e";
		when x"46" =>i:=x"5a";
		when x"47" =>i:=x"a0";
		when x"48" =>i:=x"52";
		when x"49" =>i:=x"3b";
		when x"4a" =>i:=x"d6";
		when x"4b" =>i:=x"b3";
		when x"4c" =>i:=x"29";
		when x"4d" =>i:=x"e3";
		when x"4e" =>i:=x"2f";
		when x"4f" =>i:=x"84";
		when x"50" =>i:=x"53";
		when x"51" =>i:=x"d1";
		when x"52" =>i:=x"00";
		when x"53" =>i:=x"ed";
		when x"54" =>i:=x"20";
		when x"55" =>i:=x"fc";
		when x"56" =>i:=x"b1";
		when x"57" =>i:=x"5b";
		when x"58" =>i:=x"6a";
		when x"59" =>i:=x"cb";
		when x"5a" =>i:=x"be";
		when x"5b" =>i:=x"39";
		when x"5c" =>i:=x"4a";
		when x"5d" =>i:=x"4c";
		when x"5e" =>i:=x"58";
		when x"5f" =>i:=x"cf";
		when x"60" =>i:=x"d0";
		when x"61" =>i:=x"ef";
		when x"62" =>i:=x"aa";
		when x"63" =>i:=x"fb";
		when x"64" =>i:=x"43";
		when x"65" =>i:=x"4d";
		when x"66" =>i:=x"33";
		when x"67" =>i:=x"85";
		when x"68" =>i:=x"45";
		when x"69" =>i:=x"f9";
		when x"6a" =>i:=x"02";
		when x"6b" =>i:=x"7f";
		when x"6c" =>i:=x"50";
		when x"6d" =>i:=x"3c";
		when x"6e" =>i:=x"9f";
		when x"6f" =>i:=x"a8";
		when x"70" =>i:=x"51";
		when x"71" =>i:=x"a3";
		when x"72" =>i:=x"40";
		when x"73" =>i:=x"8f";
		when x"74" =>i:=x"92";
		when x"75" =>i:=x"9d";
		when x"76" =>i:=x"38";
		when x"77" =>i:=x"f5";
		when x"78" =>i:=x"bc";
		when x"79" =>i:=x"b6";
		when x"7a" =>i:=x"da";
		when x"7b" =>i:=x"21";
		when x"7c" =>i:=x"10";
		when x"7d" =>i:=x"ff";
		when x"7e" =>i:=x"f3";
		when x"7f" =>i:=x"d2";
		when x"80" =>i:=x"cd";
		when x"81" =>i:=x"0c";
		when x"82" =>i:=x"13";
		when x"83" =>i:=x"ec";
		when x"84" =>i:=x"5f";
		when x"85" =>i:=x"97";
		when x"86" =>i:=x"44";
		when x"87" =>i:=x"17";
		when x"88" =>i:=x"c4";
		when x"89" =>i:=x"a7";
		when x"8a" =>i:=x"7e";
		when x"8b" =>i:=x"3d";
		when x"8c" =>i:=x"64";
		when x"8d" =>i:=x"5d";
		when x"8e" =>i:=x"19";
		when x"8f" =>i:=x"73";
		when x"90" =>i:=x"60";
		when x"91" =>i:=x"81";
		when x"92" =>i:=x"4f";
		when x"93" =>i:=x"dc";
		when x"94" =>i:=x"22";
		when x"95" =>i:=x"2a";
		when x"96" =>i:=x"90";
		when x"97" =>i:=x"88";
		when x"98" =>i:=x"46";
		when x"99" =>i:=x"ee";
		when x"9a" =>i:=x"b8";
		when x"9b" =>i:=x"14";
		when x"9c" =>i:=x"de";
		when x"9d" =>i:=x"5e";
		when x"9e" =>i:=x"0b";
		when x"9f" =>i:=x"db";
		when x"a0" =>i:=x"e0";
		when x"a1" =>i:=x"32";
		when x"a2" =>i:=x"3a";
		when x"a3" =>i:=x"0a";
		when x"a4" =>i:=x"49";
		when x"a5" =>i:=x"06";
		when x"a6" =>i:=x"24";
		when x"a7" =>i:=x"5c";
		when x"a8" =>i:=x"c2";
		when x"a9" =>i:=x"d3";
		when x"aa" =>i:=x"ac";
		when x"ab" =>i:=x"62";
		when x"ac" =>i:=x"91";
		when x"ad" =>i:=x"95";
		when x"ae" =>i:=x"e4";
		when x"af" =>i:=x"79";
		when x"b0" =>i:=x"e7";
		when x"b1" =>i:=x"c8";
		when x"b2" =>i:=x"37";
		when x"b3" =>i:=x"6d";
		when x"b4" =>i:=x"8d";
		when x"b5" =>i:=x"d5";
		when x"b6" =>i:=x"4e";
		when x"b7" =>i:=x"a9";
		when x"b8" =>i:=x"6c";
		when x"b9" =>i:=x"56";
		when x"ba" =>i:=x"f4";
		when x"bb" =>i:=x"ea";
		when x"bc" =>i:=x"65";
		when x"bd" =>i:=x"7a";
		when x"be" =>i:=x"ae";
		when x"bf" =>i:=x"08";
		when x"c0" =>i:=x"ba";
		when x"c1" =>i:=x"78";
		when x"c2" =>i:=x"25";
		when x"c3" =>i:=x"2e";
		when x"c4" =>i:=x"1c";
		when x"c5" =>i:=x"a6";
		when x"c6" =>i:=x"b4";
		when x"c7" =>i:=x"c6";
		when x"c8" =>i:=x"e8";
		when x"c9" =>i:=x"dd";
		when x"ca" =>i:=x"74";
		when x"cb" =>i:=x"1f";
		when x"cc" =>i:=x"4b";
		when x"cd" =>i:=x"bd";
		when x"ce" =>i:=x"8b";
		when x"cf" =>i:=x"8a";
		when x"d0" =>i:=x"70";
		when x"d1" =>i:=x"3e";
		when x"d2" =>i:=x"b5";
		when x"d3" =>i:=x"66";
		when x"d4" =>i:=x"48";
		when x"d5" =>i:=x"03";
		when x"d6" =>i:=x"f6";
		when x"d7" =>i:=x"0e";
		when x"d8" =>i:=x"61";
		when x"d9" =>i:=x"35";
		when x"da" =>i:=x"57";
		when x"db" =>i:=x"b9";
		when x"dc" =>i:=x"86";
		when x"dd" =>i:=x"c1";
		when x"de" =>i:=x"1d";
		when x"df" =>i:=x"9e";
		when x"e0" =>i:=x"e1";
		when x"e1" =>i:=x"f8";
		when x"e2" =>i:=x"98";
		when x"e3" =>i:=x"11";
		when x"e4" =>i:=x"69";
		when x"e5" =>i:=x"d9";
		when x"e6" =>i:=x"8e";
		when x"e7" =>i:=x"94";
		when x"e8" =>i:=x"9b";
		when x"e9" =>i:=x"1e";
		when x"ea" =>i:=x"87";
		when x"eb" =>i:=x"e9";
		when x"ec" =>i:=x"ce";
		when x"ed" =>i:=x"55";
		when x"ee" =>i:=x"28";
		when x"ef" =>i:=x"df";
		when x"f0" =>i:=x"8c";
		when x"f1" =>i:=x"a1";
		when x"f2" =>i:=x"89";
		when x"f3" =>i:=x"0d";
		when x"f4" =>i:=x"bf";
		when x"f5" =>i:=x"e6";
		when x"f6" =>i:=x"42";
		when x"f7" =>i:=x"68";
		when x"f8" =>i:=x"41";
		when x"f9" =>i:=x"99";
		when x"fa" =>i:=x"2d";
		when x"fb" =>i:=x"0f";
		when x"fc" =>i:=x"b0";
		when x"fd" =>i:=x"54";
		when x"fe" =>i:=x"bb";
		when x"ff" =>i:=x"16";
        when others=>null;
    end case;
    return i;
end function;
end package body util_package;
