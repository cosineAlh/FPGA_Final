--------------------------------------------

-- sbox

--------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sbox is
	Port(
		INPUT_BYTE: in STD_LOGIC_VECTOR(7 downto 0);
		OUTPUT_BYTE: out STD_LOGIC_VECTOR(7 downto 0)
	);
end sbox;

architecture Behavioral of sbox is
begin
	lut: process(INPUT_BYTE)is
	begin
		case INPUT_BYTE is
			when x"00" => OUTPUT_BYTE <= x"63";
			when x"01" => OUTPUT_BYTE <= x"7c";
			when x"02" => OUTPUT_BYTE <= x"77";
			when x"03" => OUTPUT_BYTE <= x"7b";
			when x"04" => OUTPUT_BYTE <= x"f2";
			when x"05" => OUTPUT_BYTE <= x"6b";
			when x"06" => OUTPUT_BYTE <= x"6f";
			when x"07" => OUTPUT_BYTE <= x"c5";
			when x"08" => OUTPUT_BYTE <= x"30";
			when x"09" => OUTPUT_BYTE <= x"01";
			when x"0a" => OUTPUT_BYTE <= x"67";
			when x"0b" => OUTPUT_BYTE <= x"2b";
			when x"0c" => OUTPUT_BYTE <= x"fe";
			when x"0d" => OUTPUT_BYTE <= x"d7";
			when x"0e" => OUTPUT_BYTE <= x"ab";
			when x"0f" => OUTPUT_BYTE <= x"76";
			when x"10" => OUTPUT_BYTE <= x"ca";
			when x"11" => OUTPUT_BYTE <= x"82";
			when x"12" => OUTPUT_BYTE <= x"c9";
			when x"13" => OUTPUT_BYTE <= x"7d";
			when x"14" => OUTPUT_BYTE <= x"fa";
			when x"15" => OUTPUT_BYTE <= x"59";
			when x"16" => OUTPUT_BYTE <= x"47";
			when x"17" => OUTPUT_BYTE <= x"f0";
			when x"18" => OUTPUT_BYTE <= x"ad";
			when x"19" => OUTPUT_BYTE <= x"d4";
			when x"1a" => OUTPUT_BYTE <= x"a2";
			when x"1b" => OUTPUT_BYTE <= x"af";
			when x"1c" => OUTPUT_BYTE <= x"9c";
			when x"1d" => OUTPUT_BYTE <= x"a4";
			when x"1e" => OUTPUT_BYTE <= x"72";
			when x"1f" => OUTPUT_BYTE <= x"c0";
			when x"20" => OUTPUT_BYTE <= x"b7";
			when x"21" => OUTPUT_BYTE <= x"fd";
			when x"22" => OUTPUT_BYTE <= x"93";
			when x"23" => OUTPUT_BYTE <= x"26";
			when x"24" => OUTPUT_BYTE <= x"36";
			when x"25" => OUTPUT_BYTE <= x"3f";
			when x"26" => OUTPUT_BYTE <= x"f7";
			when x"27" => OUTPUT_BYTE <= x"cc";
			when x"28" => OUTPUT_BYTE <= x"34";
			when x"29" => OUTPUT_BYTE <= x"a5";
			when x"2a" => OUTPUT_BYTE <= x"e5";
			when x"2b" => OUTPUT_BYTE <= x"f1";
			when x"2c" => OUTPUT_BYTE <= x"71";
			when x"2d" => OUTPUT_BYTE <= x"d8";
			when x"2e" => OUTPUT_BYTE <= x"31";
			when x"2f" => OUTPUT_BYTE <= x"15";
			when x"30" => OUTPUT_BYTE <= x"04";
			when x"31" => OUTPUT_BYTE <= x"c7";
			when x"32" => OUTPUT_BYTE <= x"23";
			when x"33" => OUTPUT_BYTE <= x"c3";
			when x"34" => OUTPUT_BYTE <= x"18";
			when x"35" => OUTPUT_BYTE <= x"96";
			when x"36" => OUTPUT_BYTE <= x"05";
			when x"37" => OUTPUT_BYTE <= x"9a";
			when x"38" => OUTPUT_BYTE <= x"07";
			when x"39" => OUTPUT_BYTE <= x"12";
			when x"3a" => OUTPUT_BYTE <= x"80";
			when x"3b" => OUTPUT_BYTE <= x"e2";
			when x"3c" => OUTPUT_BYTE <= x"eb";
			when x"3d" => OUTPUT_BYTE <= x"27";
			when x"3e" => OUTPUT_BYTE <= x"b2";
			when x"3f" => OUTPUT_BYTE <= x"75";
			when x"40" => OUTPUT_BYTE <= x"09";
			when x"41" => OUTPUT_BYTE <= x"83";
			when x"42" => OUTPUT_BYTE <= x"2c";
			when x"43" => OUTPUT_BYTE <= x"1a";
			when x"44" => OUTPUT_BYTE <= x"1b";
			when x"45" => OUTPUT_BYTE <= x"6e";
			when x"46" => OUTPUT_BYTE <= x"5a";
			when x"47" => OUTPUT_BYTE <= x"a0";
			when x"48" => OUTPUT_BYTE <= x"52";
			when x"49" => OUTPUT_BYTE <= x"3b";
			when x"4a" => OUTPUT_BYTE <= x"d6";
			when x"4b" => OUTPUT_BYTE <= x"b3";
			when x"4c" => OUTPUT_BYTE <= x"29";
			when x"4d" => OUTPUT_BYTE <= x"e3";
			when x"4e" => OUTPUT_BYTE <= x"2f";
			when x"4f" => OUTPUT_BYTE <= x"84";
			when x"50" => OUTPUT_BYTE <= x"53";
			when x"51" => OUTPUT_BYTE <= x"d1";
			when x"52" => OUTPUT_BYTE <= x"00";
			when x"53" => OUTPUT_BYTE <= x"ed";
			when x"54" => OUTPUT_BYTE <= x"20";
			when x"55" => OUTPUT_BYTE <= x"fc";
			when x"56" => OUTPUT_BYTE <= x"b1";
			when x"57" => OUTPUT_BYTE <= x"5b";
			when x"58" => OUTPUT_BYTE <= x"6a";
			when x"59" => OUTPUT_BYTE <= x"cb";
			when x"5a" => OUTPUT_BYTE <= x"be";
			when x"5b" => OUTPUT_BYTE <= x"39";
			when x"5c" => OUTPUT_BYTE <= x"4a";
			when x"5d" => OUTPUT_BYTE <= x"4c";
			when x"5e" => OUTPUT_BYTE <= x"58";
			when x"5f" => OUTPUT_BYTE <= x"cf";
			when x"60" => OUTPUT_BYTE <= x"d0";
			when x"61" => OUTPUT_BYTE <= x"ef";
			when x"62" => OUTPUT_BYTE <= x"aa";
			when x"63" => OUTPUT_BYTE <= x"fb";
			when x"64" => OUTPUT_BYTE <= x"43";
			when x"65" => OUTPUT_BYTE <= x"4d";
			when x"66" => OUTPUT_BYTE <= x"33";
			when x"67" => OUTPUT_BYTE <= x"85";
			when x"68" => OUTPUT_BYTE <= x"45";
			when x"69" => OUTPUT_BYTE <= x"f9";
			when x"6a" => OUTPUT_BYTE <= x"02";
			when x"6b" => OUTPUT_BYTE <= x"7f";
			when x"6c" => OUTPUT_BYTE <= x"50";
			when x"6d" => OUTPUT_BYTE <= x"3c";
			when x"6e" => OUTPUT_BYTE <= x"9f";
			when x"6f" => OUTPUT_BYTE <= x"a8";
			when x"70" => OUTPUT_BYTE <= x"51";
			when x"71" => OUTPUT_BYTE <= x"a3";
			when x"72" => OUTPUT_BYTE <= x"40";
			when x"73" => OUTPUT_BYTE <= x"8f";
			when x"74" => OUTPUT_BYTE <= x"92";
			when x"75" => OUTPUT_BYTE <= x"9d";
			when x"76" => OUTPUT_BYTE <= x"38";
			when x"77" => OUTPUT_BYTE <= x"f5";
			when x"78" => OUTPUT_BYTE <= x"bc";
			when x"79" => OUTPUT_BYTE <= x"b6";
			when x"7a" => OUTPUT_BYTE <= x"da";
			when x"7b" => OUTPUT_BYTE <= x"21";
			when x"7c" => OUTPUT_BYTE <= x"10";
			when x"7d" => OUTPUT_BYTE <= x"ff";
			when x"7e" => OUTPUT_BYTE <= x"f3";
			when x"7f" => OUTPUT_BYTE <= x"d2";
			when x"80" => OUTPUT_BYTE <= x"cd";
			when x"81" => OUTPUT_BYTE <= x"0c";
			when x"82" => OUTPUT_BYTE <= x"13";
			when x"83" => OUTPUT_BYTE <= x"ec";
			when x"84" => OUTPUT_BYTE <= x"5f";
			when x"85" => OUTPUT_BYTE <= x"97";
			when x"86" => OUTPUT_BYTE <= x"44";
			when x"87" => OUTPUT_BYTE <= x"17";
			when x"88" => OUTPUT_BYTE <= x"c4";
			when x"89" => OUTPUT_BYTE <= x"a7";
			when x"8a" => OUTPUT_BYTE <= x"7e";
			when x"8b" => OUTPUT_BYTE <= x"3d";
			when x"8c" => OUTPUT_BYTE <= x"64";
			when x"8d" => OUTPUT_BYTE <= x"5d";
			when x"8e" => OUTPUT_BYTE <= x"19";
			when x"8f" => OUTPUT_BYTE <= x"73";
			when x"90" => OUTPUT_BYTE <= x"60";
			when x"91" => OUTPUT_BYTE <= x"81";
			when x"92" => OUTPUT_BYTE <= x"4f";
			when x"93" => OUTPUT_BYTE <= x"dc";
			when x"94" => OUTPUT_BYTE <= x"22";
			when x"95" => OUTPUT_BYTE <= x"2a";
			when x"96" => OUTPUT_BYTE <= x"90";
			when x"97" => OUTPUT_BYTE <= x"88";
			when x"98" => OUTPUT_BYTE <= x"46";
			when x"99" => OUTPUT_BYTE <= x"ee";
			when x"9a" => OUTPUT_BYTE <= x"b8";
			when x"9b" => OUTPUT_BYTE <= x"14";
			when x"9c" => OUTPUT_BYTE <= x"de";
			when x"9d" => OUTPUT_BYTE <= x"5e";
			when x"9e" => OUTPUT_BYTE <= x"0b";
			when x"9f" => OUTPUT_BYTE <= x"db";
			when x"a0" => OUTPUT_BYTE <= x"e0";
			when x"a1" => OUTPUT_BYTE <= x"32";
			when x"a2" => OUTPUT_BYTE <= x"3a";
			when x"a3" => OUTPUT_BYTE <= x"0a";
			when x"a4" => OUTPUT_BYTE <= x"49";
			when x"a5" => OUTPUT_BYTE <= x"06";
			when x"a6" => OUTPUT_BYTE <= x"24";
			when x"a7" => OUTPUT_BYTE <= x"5c";
			when x"a8" => OUTPUT_BYTE <= x"c2";
			when x"a9" => OUTPUT_BYTE <= x"d3";
			when x"aa" => OUTPUT_BYTE <= x"ac";
			when x"ab" => OUTPUT_BYTE <= x"62";
			when x"ac" => OUTPUT_BYTE <= x"91";
			when x"ad" => OUTPUT_BYTE <= x"95";
			when x"ae" => OUTPUT_BYTE <= x"e4";
			when x"af" => OUTPUT_BYTE <= x"79";
			when x"b0" => OUTPUT_BYTE <= x"e7";
			when x"b1" => OUTPUT_BYTE <= x"c8";
			when x"b2" => OUTPUT_BYTE <= x"37";
			when x"b3" => OUTPUT_BYTE <= x"6d";
			when x"b4" => OUTPUT_BYTE <= x"8d";
			when x"b5" => OUTPUT_BYTE <= x"d5";
			when x"b6" => OUTPUT_BYTE <= x"4e";
			when x"b7" => OUTPUT_BYTE <= x"a9";
			when x"b8" => OUTPUT_BYTE <= x"6c";
			when x"b9" => OUTPUT_BYTE <= x"56";
			when x"ba" => OUTPUT_BYTE <= x"f4";
			when x"bb" => OUTPUT_BYTE <= x"ea";
			when x"bc" => OUTPUT_BYTE <= x"65";
			when x"bd" => OUTPUT_BYTE <= x"7a";
			when x"be" => OUTPUT_BYTE <= x"ae";
			when x"bf" => OUTPUT_BYTE <= x"08";
			when x"c0" => OUTPUT_BYTE <= x"ba";
			when x"c1" => OUTPUT_BYTE <= x"78";
			when x"c2" => OUTPUT_BYTE <= x"25";
			when x"c3" => OUTPUT_BYTE <= x"2e";
			when x"c4" => OUTPUT_BYTE <= x"1c";
			when x"c5" => OUTPUT_BYTE <= x"a6";
			when x"c6" => OUTPUT_BYTE <= x"b4";
			when x"c7" => OUTPUT_BYTE <= x"c6";
			when x"c8" => OUTPUT_BYTE <= x"e8";
			when x"c9" => OUTPUT_BYTE <= x"dd";
			when x"ca" => OUTPUT_BYTE <= x"74";
			when x"cb" => OUTPUT_BYTE <= x"1f";
			when x"cc" => OUTPUT_BYTE <= x"4b";
			when x"cd" => OUTPUT_BYTE <= x"bd";
			when x"ce" => OUTPUT_BYTE <= x"8b";
			when x"cf" => OUTPUT_BYTE <= x"8a";
			when x"d0" => OUTPUT_BYTE <= x"70";
			when x"d1" => OUTPUT_BYTE <= x"3e";
			when x"d2" => OUTPUT_BYTE <= x"b5";
			when x"d3" => OUTPUT_BYTE <= x"66";
			when x"d4" => OUTPUT_BYTE <= x"48";
			when x"d5" => OUTPUT_BYTE <= x"03";
			when x"d6" => OUTPUT_BYTE <= x"f6";
			when x"d7" => OUTPUT_BYTE <= x"0e";
			when x"d8" => OUTPUT_BYTE <= x"61";
			when x"d9" => OUTPUT_BYTE <= x"35";
			when x"da" => OUTPUT_BYTE <= x"57";
			when x"db" => OUTPUT_BYTE <= x"b9";
			when x"dc" => OUTPUT_BYTE <= x"86";
			when x"dd" => OUTPUT_BYTE <= x"c1";
			when x"de" => OUTPUT_BYTE <= x"1d";
			when x"df" => OUTPUT_BYTE <= x"9e";
			when x"e0" => OUTPUT_BYTE <= x"e1";
			when x"e1" => OUTPUT_BYTE <= x"f8";
			when x"e2" => OUTPUT_BYTE <= x"98";
			when x"e3" => OUTPUT_BYTE <= x"11";
			when x"e4" => OUTPUT_BYTE <= x"69";
			when x"e5" => OUTPUT_BYTE <= x"d9";
			when x"e6" => OUTPUT_BYTE <= x"8e";
			when x"e7" => OUTPUT_BYTE <= x"94";
			when x"e8" => OUTPUT_BYTE <= x"9b";
			when x"e9" => OUTPUT_BYTE <= x"1e";
			when x"ea" => OUTPUT_BYTE <= x"87";
			when x"eb" => OUTPUT_BYTE <= x"e9";
			when x"ec" => OUTPUT_BYTE <= x"ce";
			when x"ed" => OUTPUT_BYTE <= x"55";
			when x"ee" => OUTPUT_BYTE <= x"28";
			when x"ef" => OUTPUT_BYTE <= x"df";
			when x"f0" => OUTPUT_BYTE <= x"8c";
			when x"f1" => OUTPUT_BYTE <= x"a1";
			when x"f2" => OUTPUT_BYTE <= x"89";
			when x"f3" => OUTPUT_BYTE <= x"0d";
			when x"f4" => OUTPUT_BYTE <= x"bf";
			when x"f5" => OUTPUT_BYTE <= x"e6";
			when x"f6" => OUTPUT_BYTE <= x"42";
			when x"f7" => OUTPUT_BYTE <= x"68";
			when x"f8" => OUTPUT_BYTE <= x"41";
			when x"f9" => OUTPUT_BYTE <= x"99";
			when x"fa" => OUTPUT_BYTE <= x"2d";
			when x"fb" => OUTPUT_BYTE <= x"0f";
			when x"fc" => OUTPUT_BYTE <= x"b0";
			when x"fd" => OUTPUT_BYTE <= x"54";
			when x"fe" => OUTPUT_BYTE <= x"bb";
			when x"ff" => OUTPUT_BYTE <= x"16";
			when others => null;
		end case;
	end process;
end Behavioral;
